`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:College Of Engineering And Management 
// Student: Snehasish Biswas 
// Create Date: 11.08.2025 22:01:37
// Design Name: RTL_8-bit Arithmatic And Logic Unit 
// Module Name: alu_8bit
// Project Name: 8-bit ALU
// Target Devices: Xilinx ZYNQ 7000+ Series 
//////////////////////////////////////////////////////////////////////////////////
module alu_8bit(
    input [7:0] A,
    input [7:0] B,
    input [3:0] alu_sel,
    output [7:0] alu_out,
    output c_out
    );
reg [7:0] ALU_Result;
wire [8:0] temp;
assign alu_out=ALU_Result;
assign temp= {1'b0,A}+{1'b0,B};
assign c_out=temp[8];
always@(*)
begin 
 case(alu_sel)
    4'b0000:
     ALU_Result = A + B ; 
        4'b0001: // Subtraction
           ALU_Result = A - B ;
        4'b0010: // Multiplication
           ALU_Result = A * B;
        4'b0011: // Division
           ALU_Result = A/B;
        4'b0100: // Logical shift left
           ALU_Result = A<<1;
         4'b0101: // Logical shift right
           ALU_Result = A>>1;
         4'b0110: // Rotate left
           ALU_Result = {A[6:0],A[7]};
         4'b0111: // Rotate right
           ALU_Result = {A[0],A[7:1]};
          4'b1000: //  Logical and 
           ALU_Result = A & B;
          4'b1001: //  Logical or
           ALU_Result = A | B;
          4'b1010: //  Logical xor 
           ALU_Result = A ^ B;
          4'b1011: //  Logical nor
           ALU_Result = ~(A | B);
          4'b1100: // Logical nand 
           ALU_Result = ~(A & B);
          4'b1101: // Logical xnor
           ALU_Result = ~(A ^ B);
          4'b1110: // Greater comparison
           ALU_Result = (A>B)?8'd1:8'd0 ;
          4'b1111: // Equal comparison   
            ALU_Result = (A==B)?8'd1:8'd0 ;
          default: ALU_Result = A + B ; 
        endcase
    end

endmodule
